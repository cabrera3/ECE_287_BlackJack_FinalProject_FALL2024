module alu(
input [7:0]input_a,
input [7:0]input_b,
input [2:0]alu_control,
output reg[7:0]result);

/* build the alu */

endmodule
