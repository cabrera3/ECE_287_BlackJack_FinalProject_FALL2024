module register(
input clk, 
input rst, 
input [7:0]in, 
input en, 
output reg [7:0]out);

/* enable (en) based register */

endmodule